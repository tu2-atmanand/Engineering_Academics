-- Write the code which sir gave